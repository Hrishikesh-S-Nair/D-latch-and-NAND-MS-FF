*D_Latch 
*two tri-state inverters and a normal CMOS inverter
*----------------------------------------------
.include modelcard.pmos
.include modelcard.nmos
.model nmos nmos level=1 vto=0.5 kp=20u
.model pmos pmos level=1 vto=-0.5 kp=10u
*---------------------------------------------
* Input signals
Vd in gnd pulse(0 1.8 0 10p 10p 1n 2n)
Vclk clk gnd pulse(0 1.8 0 5p 5p 10n 20n)
*---------------------------------------------
* Tri-state inverters
*---------------------------------------------
M1 n1 n2 vdd vdd pmos L=90n W=20.0U
M2 n1 n2 gnd gnd nmos L=90n W=10.0U
M3 n3 n4 vdd vdd pmos L=90n W=20.0U
M4 n3 n4 gnd gnd nmos L=90n W=10.0U
*---------------------------------------------
* Normal CMOS inverter
*---------------------------------------------
M5 out n5 vdd vdd pmos L=90n W=20.0U
M6 out n5 gnd gnd nmos L=90n W=10.0U
*---------------------------------------------
* Capacitances
*---------------------------------------------
C1 in gnd 1f
C2 clk gnd 1f
C3 out gnd 1f
*--------------------------------------------
* Trasient Analysis
*--------------------------------------------
.tran 0.1n 100n
.control
run
plot v(in) v(clk) v(out)
.endc
.end